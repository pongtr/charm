magic
tech scmos
timestamp 1509691263
<< nwell >>
rect 53 10 91 28
<< pwell >>
rect 58 -7 95 10
<< ntransistor >>
rect 69 0 71 4
rect 77 0 79 4
<< ptransistor >>
rect 69 16 71 22
rect 77 16 79 22
<< ndiffusion >>
rect 68 0 69 4
rect 71 0 77 4
rect 79 0 80 4
<< pdiffusion >>
rect 68 18 69 22
rect 64 16 69 18
rect 71 20 77 22
rect 71 16 72 20
rect 76 16 77 20
rect 79 18 80 22
rect 79 16 84 18
<< ndcontact >>
rect 64 0 68 4
rect 80 0 84 4
<< pdcontact >>
rect 64 18 68 22
rect 72 16 76 20
rect 80 18 84 22
<< psubstratepcontact >>
rect 88 0 92 4
<< nsubstratencontact >>
rect 56 16 60 20
<< polysilicon >>
rect 69 22 71 29
rect 77 22 79 58
rect 69 4 71 16
rect 77 4 79 16
rect 69 -2 71 0
rect 77 -2 79 0
<< polycontact >>
rect 76 58 80 62
rect 80 -9 84 -5
<< metal1 >>
rect 56 20 60 28
rect 64 24 92 27
rect 64 22 68 24
rect 80 22 84 24
rect 56 -3 60 16
rect 72 12 76 16
rect 72 8 84 12
rect 80 4 84 8
rect 64 -3 68 0
rect 56 -6 68 -3
rect 80 -5 84 0
rect 88 4 92 24
rect 88 -9 92 0
<< m2contact >>
rect 76 62 80 66
rect 56 28 60 32
rect 88 -13 92 -9
<< m3contact >>
rect 56 32 60 36
rect 88 -17 92 -13
<< metal3 >>
rect 55 36 61 37
rect 55 32 56 36
rect 60 32 61 36
rect 55 31 61 32
rect 87 -13 93 -12
rect 87 -17 88 -13
rect 92 -17 93 -13
rect 87 -18 93 -17
<< labels >>
rlabel polysilicon 70 28 70 28 5 in1
rlabel polysilicon 78 28 78 28 5 in2
rlabel metal1 58 -4 58 -4 2 GND!
rlabel metal1 90 25 90 25 6 Vdd!
rlabel polycontact 82 -7 82 -7 1 out
<< end >>
