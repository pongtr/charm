magic
tech scmos
timestamp 1533067988
<< nwell >>
rect 18 18 34 31
rect -36 -4 87 18
<< pwell >>
rect -30 -33 87 -7
rect 26 -38 45 -33
<< ntransistor >>
rect -19 -21 -17 -15
rect -11 -21 -9 -15
rect 5 -21 7 -15
rect 13 -21 15 -15
rect 21 -21 23 -15
rect 29 -21 31 -15
rect 37 -21 39 -15
rect 45 -21 47 -15
rect 53 -21 55 -15
rect 69 -21 71 -15
<< ptransistor >>
rect -19 3 -17 10
rect -11 3 -9 10
rect 5 3 7 10
rect 13 3 15 10
rect 21 3 23 10
rect 29 3 31 10
rect 37 3 39 10
rect 45 3 47 10
rect 53 3 55 10
rect 69 3 71 9
<< ndiffusion >>
rect -20 -21 -19 -15
rect -17 -21 -16 -15
rect -12 -21 -11 -15
rect -9 -21 -8 -15
rect 0 -17 5 -15
rect 4 -21 5 -17
rect 7 -21 13 -15
rect 15 -19 16 -15
rect 20 -19 21 -15
rect 15 -21 21 -19
rect 23 -21 29 -15
rect 31 -21 37 -15
rect 39 -17 45 -15
rect 39 -21 40 -17
rect 44 -21 45 -17
rect 47 -21 53 -15
rect 55 -19 56 -15
rect 55 -21 60 -19
rect 68 -21 69 -15
rect 71 -21 72 -15
rect 32 -28 36 -21
<< pdiffusion >>
rect 24 10 28 21
rect -20 3 -19 10
rect -17 3 -16 10
rect -12 3 -11 10
rect -9 3 -8 10
rect 0 7 5 10
rect 4 3 5 7
rect 7 6 8 10
rect 12 6 13 10
rect 7 3 13 6
rect 15 7 21 10
rect 15 3 16 7
rect 20 3 21 7
rect 23 3 29 10
rect 31 7 37 10
rect 31 3 32 7
rect 36 3 37 7
rect 39 7 45 10
rect 39 3 40 7
rect 44 3 45 7
rect 47 6 48 10
rect 52 6 53 10
rect 47 3 53 6
rect 55 7 60 10
rect 55 3 56 7
rect 68 3 69 9
rect 71 3 72 9
<< ndcontact >>
rect -24 -21 -20 -15
rect -16 -21 -12 -15
rect -8 -21 -4 -15
rect 0 -21 4 -17
rect 16 -19 20 -15
rect 40 -21 44 -17
rect 56 -19 60 -15
rect 64 -21 68 -15
rect 72 -21 76 -15
rect 32 -32 36 -28
<< pdcontact >>
rect 24 21 28 25
rect -24 3 -20 10
rect -16 3 -12 10
rect -8 3 -4 10
rect 0 3 4 7
rect 8 6 12 10
rect 16 3 20 7
rect 32 3 36 7
rect 40 3 44 7
rect 48 6 52 10
rect 56 3 60 7
rect 64 3 68 9
rect 72 3 76 9
<< psubstratepcontact >>
rect 80 -19 84 -15
<< nsubstratencontact >>
rect -32 4 -28 8
<< polysilicon >>
rect -36 21 15 23
rect -36 15 -4 17
rect -19 10 -17 12
rect -11 10 -9 15
rect 0 17 4 18
rect 0 14 7 17
rect 5 10 7 14
rect 13 10 15 21
rect 21 10 23 12
rect 29 10 31 38
rect 37 10 39 12
rect 45 10 47 31
rect 53 21 87 23
rect 71 14 75 18
rect 79 15 87 17
rect 53 10 55 12
rect 69 9 71 11
rect -19 -15 -17 3
rect -11 -15 -9 3
rect 5 -15 7 3
rect 13 -15 15 3
rect 21 -15 23 3
rect 29 -15 31 3
rect 37 -15 39 3
rect 45 -15 47 3
rect 53 -4 55 3
rect 54 -8 55 -4
rect 53 -15 55 -8
rect 69 -15 71 3
rect -19 -35 -17 -21
rect -11 -23 -9 -21
rect 5 -23 7 -21
rect 13 -23 15 -21
rect 21 -28 23 -21
rect 29 -23 31 -21
rect 37 -35 39 -21
rect 45 -23 47 -21
rect 53 -23 55 -21
rect 69 -23 71 -21
rect -36 -37 87 -35
<< polycontact >>
rect 28 38 32 42
rect 25 31 29 35
rect -4 14 0 18
rect 44 31 48 35
rect 31 17 35 21
rect 53 17 57 21
rect 75 14 79 18
rect 50 -8 54 -4
rect 65 -8 69 -4
rect 19 -32 23 -28
<< metal1 >>
rect 32 38 43 42
rect -36 31 25 35
rect 48 31 87 35
rect -36 25 80 28
rect -36 24 24 25
rect -16 10 -12 24
rect 28 24 80 25
rect 84 24 87 28
rect 35 17 53 21
rect 8 11 52 14
rect 8 10 12 11
rect -32 -38 -28 4
rect -24 -15 -20 3
rect -8 -4 -4 3
rect 48 10 52 11
rect 0 2 4 3
rect 16 2 20 3
rect 32 2 36 3
rect 0 -1 36 2
rect 64 9 68 24
rect 40 2 44 3
rect 56 2 60 3
rect 40 -1 60 2
rect 57 -4 60 -1
rect -8 -8 50 -4
rect 57 -8 65 -4
rect -8 -15 -4 -8
rect 57 -11 60 -8
rect -24 -28 -20 -21
rect 16 -14 60 -11
rect 16 -15 20 -14
rect 56 -15 60 -14
rect 72 -15 76 3
rect 0 -22 4 -21
rect 40 -22 44 -21
rect 0 -25 44 -22
rect -24 -31 19 -28
rect -1 -32 19 -31
rect 32 -38 36 -32
rect 64 -38 68 -21
rect -36 -42 87 -38
<< m2contact >>
rect 43 38 47 42
rect 80 24 84 28
rect 0 14 4 18
rect 71 14 75 18
rect -16 -25 -12 -21
rect -16 -38 -12 -34
rect 80 -15 84 -11
rect 72 -25 76 -21
<< metal2 >>
rect 53 18 57 21
rect 4 14 71 18
rect 80 -11 84 24
rect 80 -19 84 -15
rect -16 -34 -12 -25
rect 72 -44 76 -25
<< m3contact >>
rect 47 38 51 42
<< metal3 >>
rect 46 42 52 43
rect 46 38 47 42
rect 51 38 52 42
rect 46 37 52 38
<< labels >>
rlabel polysilicon -25 -36 -25 -36 2 s
rlabel polysilicon -25 16 -25 16 3 u
rlabel polysilicon 30 34 30 34 5 a
rlabel metal1 -25 -40 -25 -40 2 GND!
rlabel metal1 -25 26 -25 26 3 Vdd!
rlabel metal2 74 -43 74 -43 8 o
rlabel metal1 4 -30 4 -30 1 _s
rlabel metal1 -2 -6 -2 -6 1 _u
rlabel polysilicon -25 22 -25 22 3 au
rlabel metal1 77 33 77 33 6 ad
rlabel metal1 -36 31 -32 35 3 ad_prev
rlabel polysilicon 85 21 87 23 7 au_next
rlabel polysilicon 85 15 87 17 7 u_next
<< end >>
