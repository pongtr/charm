magic
tech scmos
timestamp 1525658268
<< ntransistor >>
rect -43 -45 -41 -36
rect 64 -51 66 -43
rect -21 -73 -19 -61
rect -16 -73 -14 -61
rect -8 -73 -6 -61
rect -3 -73 -1 -61
rect 5 -73 7 -61
rect 13 -73 15 -61
rect 21 -73 23 -61
rect 26 -73 28 -61
rect 34 -73 36 -61
rect 39 -73 41 -61
rect -48 -83 -46 -76
<< ptransistor >>
rect -43 -24 -41 -12
rect -27 -24 -25 -12
rect -19 -24 -17 -12
rect -11 -24 -9 -12
rect -3 -24 -1 -12
rect 5 -24 7 -12
rect 13 -24 15 -12
rect 21 -24 23 -12
rect 29 -24 31 -12
rect 37 -24 39 -12
rect 45 -24 47 -12
rect 64 -24 66 -12
rect -48 -64 -46 -57
<< ndiffusion >>
rect -44 -45 -43 -36
rect -41 -45 -40 -36
rect 63 -51 64 -43
rect 66 -51 67 -43
rect -23 -66 -21 -61
rect -27 -73 -21 -66
rect -19 -73 -16 -61
rect -14 -69 -8 -61
rect -14 -73 -13 -69
rect -9 -73 -8 -69
rect -6 -73 -3 -61
rect -1 -73 0 -61
rect 4 -73 5 -61
rect 7 -73 8 -61
rect 12 -73 13 -61
rect 15 -73 16 -61
rect 20 -73 21 -61
rect 23 -73 26 -61
rect 28 -69 34 -61
rect 28 -73 29 -69
rect 33 -73 34 -69
rect 36 -73 39 -61
rect 41 -65 42 -61
rect 41 -73 46 -65
rect -49 -83 -48 -76
rect -46 -83 -45 -76
<< pdiffusion >>
rect -44 -24 -43 -12
rect -41 -24 -40 -12
rect -28 -24 -27 -12
rect -25 -24 -24 -12
rect -20 -24 -19 -12
rect -17 -24 -16 -12
rect -12 -24 -11 -12
rect -9 -16 -8 -12
rect -4 -16 -3 -12
rect -9 -24 -3 -16
rect -1 -24 0 -12
rect 4 -24 5 -12
rect 7 -24 8 -12
rect 12 -24 13 -12
rect 15 -24 16 -12
rect 20 -24 21 -12
rect 23 -16 24 -12
rect 28 -16 29 -12
rect 23 -24 29 -16
rect 31 -24 32 -12
rect 36 -24 37 -12
rect 39 -24 40 -12
rect 44 -24 45 -12
rect 47 -24 48 -12
rect 63 -24 64 -12
rect 66 -24 67 -12
rect -51 -64 -48 -57
rect -46 -64 -45 -57
<< ndcontact >>
rect -48 -45 -44 -36
rect -40 -45 -36 -36
rect 59 -51 63 -43
rect 67 -51 71 -43
rect -27 -66 -23 -61
rect -13 -73 -9 -69
rect 0 -73 4 -61
rect 8 -73 12 -61
rect 16 -73 20 -61
rect 29 -73 33 -69
rect 42 -65 46 -61
rect -53 -83 -49 -76
rect -45 -83 -41 -76
<< pdcontact >>
rect -48 -24 -44 -12
rect -40 -24 -36 -12
rect -32 -24 -28 -12
rect -24 -24 -20 -12
rect -16 -24 -12 -12
rect -8 -16 -4 -12
rect 0 -24 4 -12
rect 8 -24 12 -12
rect 16 -24 20 -12
rect 24 -16 28 -12
rect 32 -24 36 -12
rect 40 -24 44 -12
rect 48 -24 52 -12
rect 59 -24 63 -12
rect 67 -24 71 -12
rect -55 -64 -51 -57
rect -45 -64 -41 -57
<< polysilicon >>
rect -43 -12 -41 -10
rect -27 -12 -25 -10
rect -19 -12 -17 -9
rect -11 -12 -9 -10
rect -3 -12 -1 -10
rect 5 -12 7 -10
rect 13 -12 15 -10
rect 21 -12 23 -10
rect 29 -12 31 -10
rect 37 -12 39 -10
rect 45 -12 47 -10
rect 64 -12 66 -10
rect -43 -26 -41 -24
rect -27 -26 -25 -24
rect -19 -26 -17 -24
rect -11 -26 -9 -24
rect -3 -26 -1 -24
rect 5 -26 7 -24
rect 13 -26 15 -24
rect 21 -26 23 -24
rect 29 -26 31 -24
rect 37 -26 39 -24
rect 45 -26 47 -24
rect 64 -26 66 -24
rect -61 -30 -58 -28
rect -43 -36 -41 -34
rect 64 -43 66 -41
rect -43 -47 -41 -45
rect 64 -53 66 -51
rect -48 -57 -46 -55
rect -21 -61 -19 -59
rect -16 -61 -14 -59
rect -8 -61 -6 -59
rect -3 -61 -1 -59
rect 5 -61 7 -59
rect 13 -61 15 -59
rect 21 -61 23 -59
rect 26 -61 28 -59
rect 34 -61 36 -59
rect 39 -61 41 -59
rect -48 -66 -46 -64
rect -61 -71 -59 -69
rect -48 -76 -46 -74
rect -21 -75 -19 -73
rect -16 -75 -14 -73
rect -8 -75 -6 -73
rect -3 -75 -1 -73
rect 5 -75 7 -73
rect 13 -75 15 -73
rect 21 -75 23 -73
rect 26 -75 28 -73
rect 34 -75 36 -73
rect 39 -75 41 -73
rect -48 -85 -46 -83
rect -3 -111 -1 -109
rect 5 -111 7 -109
rect 13 -111 15 -109
rect 21 -111 23 -109
<< metal1 >>
rect -59 6 -55 11
rect 74 7 78 11
rect 76 -35 79 -31
rect -59 -111 -56 -106
rect 74 -111 78 -108
<< metal2 >>
rect 59 -51 63 -43
rect 67 -51 71 -43
<< labels >>
rlabel metal1 -57 10 -57 10 4 Vdd!
rlabel polysilicon -60 -29 -60 -29 1 a
rlabel metal1 76 9 76 9 6 GND!
rlabel polysilicon -60 -70 -60 -70 3 b
rlabel ndcontact -46 -41 -46 -41 1 GND!
rlabel ndcontact -51 -80 -51 -80 1 GND!
rlabel ndcontact -11 -71 -11 -71 1 GND!
rlabel ndcontact 31 -71 31 -71 1 GND!
rlabel metal2 61 -47 61 -47 1 GND!
rlabel metal1 76 -109 76 -109 8 GND!
rlabel metal1 78 -33 78 -33 7 f
rlabel metal2 69 -47 69 -47 1 f
rlabel pdcontact 69 -18 69 -18 1 f
rlabel ndcontact 10 -67 10 -67 1 _f
rlabel pdcontact 26 -14 26 -14 1 _f
rlabel pdcontact 50 -18 50 -18 1 _f
rlabel polysilicon 65 -25 65 -25 1 _f
rlabel polysilicon 65 -42 65 -42 1 _f
rlabel pdcontact -46 -18 -46 -18 1 Vdd!
rlabel pdcontact -53 -61 -53 -61 1 Vdd!
rlabel metal1 -58 -109 -58 -109 2 Vdd!
rlabel pdcontact -30 -18 -30 -18 1 Vdd!
rlabel pdcontact -6 -14 -6 -14 1 Vdd!
rlabel pdcontact 61 -18 61 -18 1 Vdd!
rlabel polysilicon -42 -11 -42 -11 1 a
rlabel polysilicon 14 -60 14 -60 1 a
rlabel polysilicon 46 -11 46 -11 1 a
rlabel polysilicon -42 -35 -42 -35 1 a
rlabel ndcontact -38 -41 -38 -41 1 _a
rlabel pdcontact -38 -18 -38 -18 1 _a
rlabel polysilicon -26 -11 -26 -11 1 _a
rlabel polysilicon 6 -60 6 -60 1 _a
rlabel polysilicon -47 -56 -47 -56 1 b
rlabel polysilicon -47 -75 -47 -75 1 b
rlabel polysilicon -7 -60 -7 -60 1 b
rlabel polysilicon 35 -60 35 -60 1 b
rlabel polysilicon -18 -11 -18 -11 1 b
rlabel polysilicon 30 -11 30 -11 1 b
rlabel polysilicon -2 -110 -2 -110 1 g0
rlabel polysilicon 6 -110 6 -110 1 g1
rlabel polysilicon 14 -110 14 -110 1 g2
rlabel polysilicon 22 -110 22 -110 1 g3
rlabel polysilicon -20 -74 -20 -74 1 g0
rlabel polysilicon -2 -74 -2 -74 1 g1
rlabel polysilicon 22 -74 22 -74 1 g2
rlabel polysilicon 40 -74 40 -74 1 g3
rlabel polysilicon -2 -11 -2 -11 5 g0
rlabel polysilicon 6 -11 6 -11 5 g1
rlabel polysilicon 14 -11 14 -11 5 g2
rlabel polysilicon 22 -11 22 -11 5 g3
rlabel pdcontact -22 -18 -22 -18 1 p1
rlabel pdcontact 10 -18 10 -18 1 p1
rlabel pdcontact 42 -18 42 -18 1 p1
rlabel pdcontact -14 -18 -14 -18 1 p2
rlabel pdcontact 2 -18 2 -18 1 p2
rlabel pdcontact 18 -18 18 -18 1 p3
rlabel pdcontact 34 -18 34 -18 1 p3
rlabel ndcontact -25 -64 -25 -64 1 n1
rlabel ndcontact 2 -67 2 -67 1 n1
rlabel ndcontact 18 -67 18 -67 1 n2
rlabel ndcontact 44 -63 44 -63 1 n2
rlabel polysilicon -15 -60 -15 -60 1 _b
rlabel polysilicon -10 -11 -10 -11 1 _b
rlabel polysilicon 38 -11 38 -11 1 _b
rlabel polysilicon 27 -60 27 -60 1 _b
rlabel ndcontact -43 -80 -43 -80 1 _b
rlabel pdcontact -43 -61 -43 -61 1 _b
<< end >>
