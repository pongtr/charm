magic
tech scmos
timestamp 1533068962
<< nwell >>
rect -10 -7 78 22
<< pwell >>
rect -2 -36 86 -7
<< ntransistor >>
rect 9 -19 11 -13
rect 25 -19 27 -13
rect 33 -19 35 -13
rect 41 -19 43 -13
rect 49 -19 51 -13
rect 65 -19 67 -13
<< ptransistor >>
rect 9 -1 11 5
rect 25 -1 27 5
rect 33 -1 35 5
rect 41 -1 43 5
rect 49 -1 51 5
rect 65 -1 67 5
<< ndiffusion >>
rect 8 -19 9 -13
rect 11 -19 12 -13
rect 24 -17 25 -13
rect 20 -19 25 -17
rect 27 -15 33 -13
rect 27 -19 28 -15
rect 32 -19 33 -15
rect 35 -19 41 -13
rect 43 -15 49 -13
rect 43 -19 44 -15
rect 48 -19 49 -15
rect 51 -19 52 -13
rect 64 -19 65 -13
rect 67 -19 68 -13
rect 36 -26 40 -19
<< pdiffusion >>
rect 28 5 32 12
rect 8 -1 9 5
rect 11 -1 12 5
rect 24 1 25 5
rect 20 -1 25 1
rect 27 -1 33 5
rect 35 -1 41 5
rect 43 3 49 5
rect 43 -1 44 3
rect 48 -1 49 3
rect 51 1 52 5
rect 51 -1 56 1
rect 64 -1 65 5
rect 67 -1 68 5
<< ndcontact >>
rect 4 -19 8 -13
rect 12 -19 16 -13
rect 20 -17 24 -13
rect 28 -19 32 -15
rect 44 -19 48 -15
rect 52 -19 56 -13
rect 60 -19 64 -13
rect 68 -19 72 -13
rect 36 -30 40 -26
<< pdcontact >>
rect 28 12 32 16
rect 4 -1 8 5
rect 12 -1 16 5
rect 20 1 24 5
rect 44 -1 48 3
rect 52 1 56 5
rect 60 -1 64 5
rect 68 -1 72 5
<< psubstratepcontact >>
rect 76 -17 80 -13
<< nsubstratencontact >>
rect -4 -1 0 3
<< polysilicon >>
rect 9 9 11 22
rect 9 7 27 9
rect 9 5 11 7
rect 25 5 27 7
rect 33 5 35 7
rect 41 5 43 7
rect 49 5 51 7
rect 65 5 67 7
rect 9 -13 11 -1
rect 25 -13 27 -1
rect 33 -2 35 -1
rect 33 -13 35 -6
rect 41 -13 43 -1
rect 49 -13 51 -1
rect 65 -13 67 -1
rect 9 -21 11 -19
rect 25 -21 27 -19
rect 33 -21 35 -19
rect 41 -24 43 -19
rect 49 -21 51 -19
rect 65 -24 67 -19
rect 41 -26 67 -24
rect 41 -31 43 -26
rect -10 -33 43 -31
<< polycontact >>
rect 31 -6 35 -2
rect 51 -6 55 -2
<< metal1 >>
rect 76 16 80 22
rect 4 12 28 16
rect 32 12 80 16
rect 4 5 8 12
rect 20 6 56 9
rect 20 5 24 6
rect 52 5 56 6
rect 68 5 72 12
rect -4 -26 0 -1
rect 12 -2 16 -1
rect 12 -6 31 -2
rect 12 -13 16 -6
rect 44 -9 48 -1
rect 60 -2 64 -1
rect 55 -6 64 -2
rect 20 -12 56 -9
rect 20 -13 24 -12
rect 52 -13 56 -12
rect 4 -26 8 -19
rect 28 -22 48 -19
rect 60 -13 64 -6
rect 76 -13 80 12
rect 68 -26 72 -19
rect -4 -30 36 -26
rect 40 -30 72 -26
rect -4 -36 0 -30
<< m2contact >>
rect 52 -23 56 -19
<< metal2 >>
rect 52 -36 56 -23
<< labels >>
rlabel metal1 6 -28 6 -28 3 GND!
rlabel metal1 6 14 6 14 4 Vdd!
rlabel polysilicon 10 17 10 17 5 b
rlabel polysilicon 3 -32 3 -32 2 cin
rlabel metal2 54 -33 54 -33 1 o
<< end >>
