magic
tech scmos
timestamp 1533662855
<< nwell >>
rect 14 39 171 58
<< pwell >>
rect 7 17 166 36
<< ntransistor >>
rect 26 23 28 30
rect 35 23 37 30
rect 43 23 45 30
rect 59 23 61 30
rect 75 23 90 30
rect 104 23 106 30
rect 112 23 114 30
rect 128 23 130 30
rect 144 23 146 30
rect 152 23 154 30
<< ptransistor >>
rect 26 45 28 52
rect 35 45 37 52
rect 43 45 45 52
rect 59 45 61 52
rect 75 45 90 52
rect 104 45 106 52
rect 112 45 114 52
rect 128 45 130 52
rect 144 45 146 52
rect 152 45 154 52
<< ndiffusion >>
rect 24 23 26 30
rect 28 27 35 30
rect 28 23 30 27
rect 34 23 35 27
rect 37 26 38 30
rect 42 26 43 30
rect 37 23 43 26
rect 45 26 46 30
rect 45 23 50 26
rect 54 27 59 30
rect 58 23 59 27
rect 61 26 62 30
rect 61 23 66 26
rect 70 27 75 30
rect 74 23 75 27
rect 90 26 91 30
rect 90 23 95 26
rect 99 27 104 30
rect 103 23 104 27
rect 106 23 107 30
rect 111 23 112 30
rect 114 26 115 30
rect 114 23 119 26
rect 123 27 128 30
rect 127 23 128 27
rect 130 26 131 30
rect 130 23 135 26
rect 143 23 144 30
rect 146 27 152 30
rect 146 23 147 27
rect 151 23 152 27
rect 154 23 155 30
<< pdiffusion >>
rect 20 49 26 52
rect 24 45 26 49
rect 28 48 30 52
rect 34 48 35 52
rect 28 45 35 48
rect 37 49 43 52
rect 37 45 38 49
rect 42 45 43 49
rect 45 49 50 52
rect 45 45 46 49
rect 58 48 59 52
rect 54 45 59 48
rect 61 49 66 52
rect 61 45 62 49
rect 74 48 75 52
rect 70 45 75 48
rect 90 49 95 52
rect 90 45 91 49
rect 103 48 104 52
rect 99 45 104 48
rect 106 45 107 52
rect 111 45 112 52
rect 114 49 119 52
rect 114 45 115 49
rect 127 48 128 52
rect 123 45 128 48
rect 130 49 135 52
rect 130 45 131 49
rect 139 49 144 52
rect 143 45 144 49
rect 146 48 147 52
rect 151 48 152 52
rect 146 45 152 48
rect 154 49 159 52
rect 154 45 155 49
<< ndcontact >>
rect 20 23 24 30
rect 30 23 34 27
rect 38 26 42 30
rect 46 26 50 30
rect 54 23 58 27
rect 62 26 66 30
rect 70 23 74 27
rect 91 26 95 30
rect 99 23 103 27
rect 107 23 111 30
rect 115 26 119 30
rect 123 23 127 27
rect 131 26 135 30
rect 139 23 143 30
rect 147 23 151 27
rect 155 23 159 30
<< pdcontact >>
rect 20 45 24 49
rect 30 48 34 52
rect 38 45 42 49
rect 46 45 50 49
rect 54 48 58 52
rect 62 45 66 49
rect 70 48 74 52
rect 91 45 95 49
rect 99 48 103 52
rect 107 45 111 52
rect 115 45 119 49
rect 123 48 127 52
rect 131 45 135 49
rect 139 45 143 49
rect 147 48 151 52
rect 155 45 159 49
<< psubstratepcontact >>
rect 10 20 14 24
<< nsubstratencontact >>
rect 164 47 168 51
<< polysilicon >>
rect 26 59 28 66
rect 152 62 154 66
rect 112 60 154 62
rect 26 57 45 59
rect 26 52 28 57
rect 35 52 37 54
rect 43 52 45 57
rect 59 52 61 54
rect 75 52 90 54
rect 104 52 106 54
rect 112 52 114 60
rect 128 53 135 55
rect 139 53 146 55
rect 128 52 130 53
rect 144 52 146 53
rect 152 52 154 60
rect 26 34 28 45
rect 16 32 28 34
rect 16 9 18 32
rect 26 30 28 32
rect 35 30 37 45
rect 43 43 45 45
rect 43 30 45 32
rect 59 30 61 45
rect 75 30 90 45
rect 104 30 106 45
rect 112 43 114 45
rect 128 43 130 45
rect 112 30 114 32
rect 128 30 130 32
rect 144 30 146 45
rect 152 30 154 45
rect 26 21 28 23
rect 35 21 37 23
rect 43 18 45 23
rect 59 21 61 23
rect 75 21 90 23
rect 104 21 106 23
rect 25 16 45 18
rect 112 15 114 23
rect 128 19 130 23
rect 128 17 135 19
rect 16 7 28 9
rect 26 0 28 7
rect 144 4 146 23
rect 139 2 146 4
rect 152 0 154 23
<< polycontact >>
rect 135 53 139 57
rect 31 40 35 44
rect 55 35 59 39
rect 71 40 75 44
rect 100 31 104 35
rect 21 14 25 18
rect 135 17 139 21
rect 112 11 116 15
rect 135 0 139 4
<< metal1 >>
rect 14 64 17 66
rect 14 60 30 64
rect 14 0 17 60
rect 30 52 34 60
rect 54 52 58 60
rect 20 30 24 45
rect 38 30 42 45
rect 70 52 74 60
rect 46 39 50 45
rect 99 52 103 60
rect 135 57 139 66
rect 62 44 66 45
rect 107 52 127 55
rect 62 40 71 44
rect 46 31 55 39
rect 46 30 50 31
rect 62 30 66 40
rect 20 22 25 23
rect 21 18 25 22
rect 30 10 34 23
rect 91 35 95 45
rect 95 31 100 35
rect 91 30 95 31
rect 54 10 58 23
rect 107 30 111 45
rect 70 10 74 23
rect 99 10 103 23
rect 147 52 151 60
rect 115 44 119 45
rect 115 30 119 40
rect 131 35 135 45
rect 131 30 135 31
rect 162 51 166 66
rect 139 30 143 45
rect 107 20 127 23
rect 155 30 159 45
rect 139 17 143 23
rect 155 14 159 23
rect 116 11 159 14
rect 162 47 164 51
rect 162 10 166 47
rect 162 0 166 6
<< m2contact >>
rect 30 60 34 64
rect 54 60 58 64
rect 27 40 31 44
rect 70 60 74 64
rect 99 60 103 64
rect 147 60 151 64
rect 55 31 59 35
rect 30 6 34 10
rect 91 31 95 35
rect 54 6 58 10
rect 70 6 74 10
rect 115 40 119 44
rect 131 31 135 35
rect 147 19 151 23
rect 99 6 103 10
rect 162 6 166 10
<< metal2 >>
rect 34 60 54 64
rect 58 60 70 64
rect 74 60 99 64
rect 103 60 147 64
rect 173 44 177 52
rect 1 40 27 44
rect 119 40 177 44
rect 1 39 6 40
rect 59 31 91 35
rect 135 31 177 35
rect 34 6 54 9
rect 58 6 70 9
rect 74 6 99 9
rect 147 9 151 19
rect 173 14 177 31
rect 103 6 162 9
<< m3contact >>
rect 173 52 177 56
rect 1 34 6 39
rect 173 10 177 14
<< metal3 >>
rect 172 56 178 57
rect 172 52 173 56
rect 177 52 178 56
rect 172 51 178 52
rect 0 39 7 40
rect 0 34 1 39
rect 6 34 7 39
rect 0 33 7 34
rect 172 14 178 15
rect 172 10 173 14
rect 177 10 178 14
rect 172 9 178 10
<< labels >>
rlabel polysilicon 27 65 27 65 5 w
rlabel metal1 15 65 15 65 4 Vdd!
rlabel metal2 13 42 13 42 3 in
rlabel metal2 167 33 167 33 7 port1
rlabel metal1 137 65 137 65 5 r1
rlabel polysilicon 153 65 153 65 5 r0
rlabel metal1 164 65 164 65 6 GND!
rlabel metal2 167 42 167 42 7 port0
rlabel polysilicon 26 0 28 2 1 w_next
rlabel polycontact 135 0 139 4 1 r1_next
rlabel polysilicon 152 0 154 2 1 r0_next
<< end >>
