magic
tech scmos
timestamp 1525671357
<< ntransistor >>
rect 5 0 7 3
rect 5 -10 7 -7
rect 5 -62 7 -59
rect 5 -72 7 -69
<< ptransistor >>
rect 5 15 7 21
rect 5 -29 7 -23
rect 5 -47 7 -41
rect 5 -91 7 -85
<< ndiffusion >>
rect 4 0 5 3
rect 7 0 8 3
rect 4 -10 5 -7
rect 7 -10 8 -7
rect 4 -62 5 -59
rect 7 -62 8 -59
rect 4 -72 5 -69
rect 7 -72 8 -69
<< pdiffusion >>
rect 4 17 5 21
rect 0 15 5 17
rect 7 19 12 21
rect 7 15 8 19
rect 4 -29 5 -23
rect 7 -27 8 -23
rect 7 -29 12 -27
rect 0 -43 5 -41
rect 4 -47 5 -43
rect 7 -45 8 -41
rect 7 -47 12 -45
rect 4 -89 5 -85
rect 0 -91 5 -89
rect 7 -89 8 -85
rect 7 -91 12 -89
<< ndcontact >>
rect 0 -1 4 3
rect 8 -1 12 3
rect 0 -11 4 -7
rect 8 -11 12 -7
rect 0 -63 4 -59
rect 8 -63 12 -59
rect 0 -73 4 -69
rect 8 -73 12 -69
<< pdcontact >>
rect 0 17 4 21
rect 8 15 12 19
rect 0 -29 4 -23
rect 8 -27 12 -23
rect 0 -47 4 -43
rect 8 -45 12 -41
rect 0 -89 4 -85
rect 8 -89 12 -85
<< polysilicon >>
rect 5 21 7 23
rect 5 13 7 15
rect 5 3 7 5
rect 5 -2 7 0
rect 5 -7 7 -5
rect 5 -12 7 -10
rect -9 -14 -7 -12
rect 16 -14 18 -12
rect -9 -21 -7 -19
rect 16 -21 18 -19
rect 5 -23 7 -21
rect 5 -31 7 -29
rect 5 -41 7 -39
rect 5 -49 7 -47
rect 5 -59 7 -57
rect 5 -64 7 -62
rect 5 -69 7 -67
rect 5 -74 7 -72
rect -9 -76 -6 -74
rect 16 -76 18 -74
rect -9 -83 -6 -81
rect 16 -83 18 -81
rect 5 -85 7 -83
rect 5 -93 7 -91
<< metal1 >>
rect -6 25 -3 28
rect -9 -63 -6 -59
rect 16 -63 19 -59
rect -9 -96 -3 -93
rect 15 -96 18 -93
rect -6 -98 -3 -96
<< m2contact >>
rect 15 -89 19 -85
<< metal2 >>
rect -9 22 -6 25
rect 16 22 19 25
rect -9 -89 -6 -85
<< labels >>
rlabel metal2 -9 -87 -9 -87 3 i0
rlabel metal1 -8 -95 -8 -95 2 GND!
rlabel metal2 -8 23 -8 23 4 Vdd!
rlabel polysilicon -9 -14 -9 -12 3 c0
rlabel polysilicon -9 -21 -9 -19 3 _c0
rlabel polysilicon -9 -76 -9 -74 3 c1
rlabel polysilicon -9 -83 -9 -81 3 _c1
rlabel pdcontact 2 19 2 19 1 Vdd!
rlabel metal2 17 23 17 23 6 Vdd!
rlabel metal1 -5 26 -5 26 4 GND!
rlabel metal1 17 -95 17 -95 8 GND!
rlabel metal1 18 -61 18 -61 7 GND2!
rlabel metal1 -7 -61 -7 -61 3 GND!
rlabel pdcontact 10 -25 10 -25 1 connection1
rlabel ndcontact 10 -9 10 -9 1 connection1
rlabel ndcontact 10 1 10 1 1 connection1
rlabel pdcontact 10 17 10 17 1 connection1
rlabel ndcontact 2 -9 2 -9 1 connection2
rlabel pdcontact 2 -26 2 -26 1 connection2
rlabel polysilicon 6 -40 6 -40 1 connection2
rlabel polysilicon 6 -58 6 -58 1 connection2
rlabel pdcontact 2 -45 2 -45 1 connection3
rlabel ndcontact 2 -61 2 -61 1 connection3
rlabel ndcontact 2 -71 2 -71 1 connection3
rlabel pdcontact 2 -87 2 -87 1 connection3
rlabel pdcontact 10 -43 10 -43 1 Vdd!
rlabel ndcontact 2 1 2 1 1 GND!
rlabel polysilicon 6 14 6 14 1 i0
rlabel polysilicon 6 -1 6 -1 1 i0
rlabel ndcontact 10 -71 10 -71 1 out
rlabel pdcontact 10 -87 10 -87 1 out
rlabel m2contact 17 -87 17 -87 7 out
rlabel polysilicon 6 -84 6 -84 1 _c1
rlabel polysilicon 6 -73 6 -73 1 c1
rlabel polysilicon 17 -75 17 -75 7 c1
rlabel polysilicon 17 -82 17 -82 7 _c1
rlabel polysilicon 17 -20 17 -20 7 _c0
rlabel polysilicon 6 -6 6 -6 1 c0
rlabel polysilicon 17 -13 17 -13 7 c0
rlabel ndcontact 10 -61 10 -61 1 GND2!
rlabel polysilicon 6 -22 6 -22 1 _c0
<< end >>
