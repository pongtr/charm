magic
tech scmos
timestamp 1525667722
<< error_p >>
rect -46 1251 -43 1252
<< ntransistor >>
rect -22 1296 -20 1303
rect -4 1296 -2 1303
rect 14 1296 16 1303
rect 32 1296 34 1303
rect 49 1296 51 1303
rect 68 1296 70 1303
<< ptransistor >>
rect -22 1326 -20 1333
rect -4 1326 -2 1333
rect 14 1326 16 1333
rect 32 1326 34 1333
rect 49 1326 51 1333
rect 68 1326 70 1333
<< ndiffusion >>
rect -28 1301 -22 1303
rect -23 1296 -22 1301
rect -20 1298 -19 1303
rect -20 1296 -14 1298
rect -5 1298 -4 1303
rect -10 1296 -4 1298
rect -2 1298 -1 1303
rect -2 1296 4 1298
rect 8 1301 14 1303
rect 13 1296 14 1301
rect 16 1298 17 1303
rect 16 1296 22 1298
rect 26 1301 32 1303
rect 31 1296 32 1301
rect 34 1298 35 1303
rect 40 1298 49 1303
rect 34 1296 49 1298
rect 51 1298 54 1303
rect 51 1296 59 1298
rect 67 1299 68 1303
rect 63 1296 68 1299
rect 70 1299 71 1303
rect 70 1296 75 1299
<< pdiffusion >>
rect -23 1328 -22 1333
rect -28 1326 -22 1328
rect -20 1331 -14 1333
rect -20 1326 -19 1331
rect -10 1331 -4 1333
rect -5 1326 -4 1331
rect -2 1331 4 1333
rect -2 1326 -1 1331
rect 13 1328 14 1333
rect 8 1326 14 1328
rect 16 1331 22 1333
rect 16 1326 17 1331
rect 31 1328 32 1333
rect 26 1326 32 1328
rect 34 1331 49 1333
rect 34 1326 35 1331
rect 40 1326 49 1331
rect 51 1331 59 1333
rect 51 1326 54 1331
rect 63 1330 68 1333
rect 67 1326 68 1330
rect 70 1330 75 1333
rect 70 1326 71 1330
<< ndcontact >>
rect -28 1296 -23 1301
rect -19 1298 -14 1303
rect -10 1298 -5 1303
rect -1 1298 4 1303
rect 8 1296 13 1301
rect 17 1298 22 1303
rect 26 1296 31 1301
rect 35 1298 40 1303
rect 54 1298 59 1303
rect 63 1299 67 1303
rect 71 1299 75 1303
<< pdcontact >>
rect -28 1328 -23 1333
rect -19 1326 -14 1331
rect -10 1326 -5 1331
rect -1 1326 4 1331
rect 8 1328 13 1333
rect 17 1326 22 1331
rect 26 1328 31 1333
rect 35 1326 40 1331
rect 54 1326 59 1331
rect 63 1326 67 1330
rect 71 1326 75 1330
<< polysilicon >>
rect -22 1333 -20 1335
rect -4 1333 -2 1335
rect 14 1333 16 1335
rect 32 1333 34 1335
rect 49 1333 51 1335
rect 68 1333 70 1335
rect -22 1324 -20 1326
rect -4 1324 -2 1326
rect 14 1324 16 1326
rect 32 1324 34 1326
rect 49 1324 51 1326
rect 68 1324 70 1326
rect -22 1303 -20 1305
rect -4 1303 -2 1305
rect 14 1303 16 1305
rect 32 1303 34 1305
rect 49 1303 51 1305
rect 68 1303 70 1306
rect -22 1294 -20 1296
rect -4 1294 -2 1296
rect 14 1294 16 1296
rect 32 1294 34 1296
rect 49 1294 51 1296
rect 68 1294 70 1296
<< metal1 >>
rect -46 1369 -43 1373
rect 82 1369 85 1373
rect 80 1327 85 1332
rect -40 1315 -35 1319
rect -46 1297 -41 1302
rect -46 1249 -43 1251
rect -35 1249 -31 1252
rect 82 1249 85 1254
<< m2contact >>
rect -35 1369 -31 1373
<< metal2 >>
rect -40 1308 -36 1312
<< labels >>
rlabel metal2 -39 1310 -39 1310 1 in
rlabel metal1 -39 1317 -39 1317 1 CLK
rlabel metal1 -43 1299 -43 1299 3 Vdd!
rlabel pdcontact -26 1330 -26 1330 1 Vdd!
rlabel pdcontact 10 1331 10 1331 1 Vdd!
rlabel pdcontact 29 1330 29 1330 1 Vdd!
rlabel metal1 -45 1372 -45 1372 4 Vdd!
rlabel metal1 -45 1250 -45 1250 2 Vdd!
rlabel ndcontact -26 1298 -26 1298 1 GND!
rlabel ndcontact 11 1298 11 1298 1 GND!
rlabel ndcontact 28 1298 28 1298 1 GND!
rlabel metal1 83 1251 83 1251 1 GND!
rlabel metal1 82 1329 82 1329 1 GND!
rlabel metal1 83 1371 83 1371 5 GND!
rlabel polysilicon -21 1334 -21 1334 1 CLK
rlabel polysilicon -21 1295 -21 1295 1 CLK
rlabel polysilicon -3 1304 -3 1304 1 CLK
rlabel polysilicon 50 1334 50 1334 1 CLK
rlabel polysilicon 69 1304 69 1304 1 CLK
rlabel m2contact -33 1371 -33 1371 5 CLK
rlabel metal1 -33 1250 -33 1250 1 CLK
rlabel ndcontact -17 1300 -17 1301 1 _CLK
rlabel pdcontact -16 1328 -16 1328 1 _CLK
rlabel polysilicon -3 1334 -3 1334 1 _CLK
rlabel polysilicon 50 1304 50 1304 1 _CLK
rlabel polysilicon 69 1334 69 1334 1 _CLK
rlabel ndcontact -7 1300 -7 1300 1 in
rlabel pdcontact -8 1329 -8 1329 1 in
rlabel pdcontact 1 1328 1 1328 1 stage1
rlabel ndcontact 1 1300 1 1300 1 stage1
rlabel polysilicon 15 1325 15 1325 1 stage1
rlabel polysilicon 15 1304 15 1304 1 stage1
rlabel ndcontact 57 1301 57 1301 1 stage1
rlabel pdcontact 57 1328 57 1328 1 stage1
rlabel pdcontact 65 1327 65 1327 1 stage1
rlabel ndcontact 65 1301 65 1301 1 stage1
rlabel pdcontact 20 1328 20 1328 1 stage2
rlabel ndcontact 20 1300 20 1300 1 stage2
rlabel pdcontact 37 1328 37 1328 1 stage2
rlabel ndcontact 37 1300 37 1300 1 stage2
rlabel pdcontact 73 1327 73 1327 1 out
rlabel ndcontact 73 1301 73 1301 1 out
<< end >>
