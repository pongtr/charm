magic
tech scmos
timestamp 1525668657
<< ntransistor >>
rect -19 -21 -17 -15
rect -11 -21 -9 -15
rect 5 -21 7 -15
rect 13 -21 15 -15
rect 21 -21 23 -15
rect 29 -21 31 -15
rect 37 -21 39 -15
rect 45 -21 47 -15
rect 53 -21 55 -15
rect 69 -21 71 -15
<< ptransistor >>
rect -19 3 -17 10
rect -11 3 -9 10
rect 5 3 7 10
rect 13 3 15 10
rect 21 3 23 10
rect 29 3 31 10
rect 37 3 39 10
rect 45 3 47 10
rect 53 3 55 10
rect 69 3 71 9
<< ndiffusion >>
rect -20 -21 -19 -15
rect -17 -21 -16 -15
rect -12 -21 -11 -15
rect -9 -21 -8 -15
rect 0 -17 5 -15
rect 4 -21 5 -17
rect 7 -21 13 -15
rect 15 -19 16 -15
rect 20 -19 21 -15
rect 15 -21 21 -19
rect 23 -21 29 -15
rect 31 -21 37 -15
rect 39 -17 45 -15
rect 39 -21 40 -17
rect 44 -21 45 -17
rect 47 -21 53 -15
rect 55 -19 56 -15
rect 55 -21 60 -19
rect 68 -21 69 -15
rect 71 -21 72 -15
rect 32 -28 36 -21
<< pdiffusion >>
rect 24 10 28 21
rect -20 3 -19 10
rect -17 3 -16 10
rect -12 3 -11 10
rect -9 3 -8 10
rect 0 7 5 10
rect 4 3 5 7
rect 7 6 8 10
rect 12 6 13 10
rect 7 3 13 6
rect 15 7 21 10
rect 15 3 16 7
rect 20 3 21 7
rect 23 3 29 10
rect 31 7 37 10
rect 31 3 32 7
rect 36 3 37 7
rect 39 7 45 10
rect 39 3 40 7
rect 44 3 45 7
rect 47 6 48 10
rect 52 6 53 10
rect 47 3 53 6
rect 55 7 60 10
rect 55 3 56 7
rect 68 3 69 9
rect 71 3 72 9
<< ndcontact >>
rect -24 -21 -20 -15
rect -16 -21 -12 -15
rect -8 -21 -4 -15
rect 0 -21 4 -17
rect 16 -19 20 -15
rect 40 -21 44 -17
rect 56 -19 60 -15
rect 64 -21 68 -15
rect 72 -21 76 -15
rect 32 -32 36 -28
<< pdcontact >>
rect 24 21 28 25
rect -24 3 -20 10
rect -16 3 -12 10
rect -8 3 -4 10
rect 0 3 4 7
rect 8 6 12 10
rect 16 3 20 7
rect 32 3 36 7
rect 40 3 44 7
rect 48 6 52 10
rect 56 3 60 7
rect 64 3 68 9
rect 72 3 76 9
<< polysilicon >>
rect -26 21 -23 23
rect 77 21 80 23
rect -26 15 -23 17
rect -19 10 -17 12
rect -11 10 -9 12
rect 5 10 7 12
rect 13 10 15 12
rect 21 10 23 12
rect 78 15 80 17
rect 29 10 31 12
rect 37 10 39 12
rect 45 10 47 12
rect 53 10 55 12
rect 69 9 71 11
rect -19 1 -17 3
rect -11 1 -9 3
rect 5 1 7 3
rect 13 1 15 3
rect 21 1 23 3
rect 29 1 31 3
rect 37 1 39 3
rect 45 1 47 3
rect 53 1 55 3
rect 69 1 71 3
rect -19 -15 -17 -13
rect -11 -15 -9 -13
rect 5 -15 7 -13
rect 13 -15 15 -13
rect 21 -15 23 -13
rect 29 -15 31 -13
rect 37 -15 39 -13
rect 45 -15 47 -13
rect 53 -15 55 -13
rect 69 -15 71 -13
rect -19 -23 -17 -21
rect -11 -23 -9 -21
rect 5 -23 7 -21
rect 13 -23 15 -21
rect 21 -23 23 -21
rect 29 -23 31 -21
rect 37 -23 39 -21
rect 45 -23 47 -21
rect 53 -23 55 -21
rect 69 -23 71 -21
rect -26 -37 -24 -35
rect 77 -37 80 -35
<< metal1 >>
rect -26 31 -23 35
rect 77 31 80 35
rect -26 24 -22 28
rect 77 24 80 28
rect -26 -42 -23 -38
rect 77 -42 80 -38
<< metal2 >>
rect 72 -44 76 -41
<< labels >>
rlabel polysilicon -25 -36 -25 -36 2 s
rlabel polysilicon -25 16 -25 16 3 u
rlabel metal1 -25 -40 -25 -40 2 GND!
rlabel metal1 -25 26 -25 26 3 Vdd!
rlabel metal2 74 -43 74 -43 8 o
rlabel polysilicon -25 22 -25 22 3 au
rlabel pdcontact -14 6 -14 6 1 Vdd!
rlabel pdcontact 26 23 26 23 1 Vdd!
rlabel pdcontact 66 6 66 6 1 Vdd!
rlabel metal1 78 26 78 26 7 Vdd!
rlabel ndcontact -14 -18 -14 -18 1 GND!
rlabel ndcontact 34 -30 34 -30 1 GND!
rlabel ndcontact 66 -18 66 -18 1 GND!
rlabel metal1 79 -40 79 -40 8 GND!
rlabel polysilicon -18 -14 -18 -14 1 s
rlabel polysilicon -18 11 -18 11 1 s
rlabel polysilicon -10 11 -10 11 1 u
rlabel polysilicon -10 -14 -10 -14 1 u
rlabel ndcontact 2 -19 2 -19 1 n1
rlabel ndcontact 42 -19 42 -19 1 n1
rlabel pdcontact 2 5 2 5 1 p1
rlabel pdcontact 18 5 18 5 1 p1
rlabel pdcontact 34 5 34 5 1 p1
rlabel pdcontact 10 8 10 8 1 p2
rlabel pdcontact 50 8 50 8 1 p2
rlabel ndcontact -6 -18 -6 -18 1 _u
rlabel pdcontact -6 7 -6 7 1 _u
rlabel polysilicon 54 -22 54 -22 1 _u
rlabel polysilicon 54 11 54 11 1 _u
rlabel polysilicon 6 11 6 11 1 u
rlabel polysilicon 6 -14 6 -14 1 u
rlabel polysilicon 79 16 79 16 7 u
rlabel pdcontact -22 6 -22 6 3 _s
rlabel ndcontact -22 -18 -22 -18 3 _s
rlabel polysilicon 22 -22 22 -22 1 _s
rlabel polysilicon 22 11 22 11 1 _s
rlabel polysilicon 14 -14 14 -14 1 au
rlabel polysilicon 14 11 14 11 1 au
rlabel ndcontact 18 -17 18 -17 1 _o
rlabel ndcontact 58 -17 58 -17 1 _o
rlabel pdcontact 42 5 42 5 1 _o
rlabel pdcontact 58 5 58 5 1 _o
rlabel polysilicon 70 -14 70 -14 1 _o
rlabel polysilicon 70 2 70 2 1 _o
rlabel pdcontact 74 6 74 6 1 o
rlabel ndcontact 74 -18 74 -18 1 o
rlabel polysilicon 79 -36 79 -36 7 s
rlabel polysilicon 38 11 38 11 1 s
rlabel polysilicon 38 -22 38 -22 1 s
rlabel polysilicon 46 -22 46 -22 1 ad
rlabel polysilicon 46 11 46 11 1 ad
rlabel polysilicon 30 11 30 11 1 a
rlabel polysilicon 30 -14 30 -14 1 a
rlabel metal1 -25 33 -25 33 4 a
rlabel polysilicon 79 22 79 22 7 a
rlabel metal1 78 33 78 33 6 ad
<< end >>
