magic
tech scmos
timestamp 1533067988
<< nwell >>
rect -58 -30 85 -6
rect -69 -70 -35 -51
<< pwell >>
rect -59 -51 79 -30
rect -33 -70 77 -51
rect -59 -74 77 -70
rect -59 -99 75 -74
<< ntransistor >>
rect -43 -45 -41 -36
rect -48 -83 -46 -76
rect -21 -73 -19 -61
rect -16 -73 -14 -61
rect -8 -73 -6 -61
rect -3 -73 -1 -61
rect 5 -73 7 -61
rect 13 -73 15 -61
rect 21 -73 23 -61
rect 26 -62 31 -61
rect 26 -73 28 -62
rect 34 -73 36 -61
rect 39 -73 41 -61
rect 64 -51 66 -43
<< ptransistor >>
rect -43 -24 -41 -12
rect -27 -24 -25 -12
rect -19 -24 -17 -12
rect -11 -24 -9 -12
rect -3 -24 -1 -12
rect 5 -24 7 -12
rect 13 -24 15 -12
rect 21 -24 23 -12
rect 29 -24 31 -12
rect 37 -24 39 -12
rect 45 -24 47 -12
rect 64 -24 66 -12
rect -48 -64 -46 -57
<< ndiffusion >>
rect -44 -45 -43 -36
rect -41 -45 -40 -36
rect -49 -83 -48 -76
rect -46 -83 -45 -76
rect -23 -66 -21 -61
rect -27 -73 -21 -66
rect -19 -73 -16 -61
rect -14 -69 -8 -61
rect -14 -73 -13 -69
rect -9 -73 -8 -69
rect -6 -73 -3 -61
rect -1 -73 0 -61
rect 4 -73 5 -61
rect 7 -73 8 -61
rect 12 -73 13 -61
rect 15 -73 16 -61
rect 20 -73 21 -61
rect 23 -73 26 -61
rect 31 -62 34 -61
rect 28 -69 34 -62
rect 28 -73 29 -69
rect 33 -73 34 -69
rect 36 -73 39 -61
rect 41 -65 42 -61
rect 41 -73 46 -65
rect 63 -51 64 -43
rect 66 -51 67 -43
<< pdiffusion >>
rect -44 -24 -43 -12
rect -41 -24 -40 -12
rect -28 -24 -27 -12
rect -25 -24 -24 -12
rect -20 -24 -19 -12
rect -17 -24 -16 -12
rect -12 -24 -11 -12
rect -9 -16 -8 -12
rect -4 -16 -3 -12
rect -9 -24 -3 -16
rect -1 -24 0 -12
rect 4 -24 5 -12
rect 7 -24 8 -12
rect 12 -24 13 -12
rect 15 -24 16 -12
rect 20 -24 21 -12
rect 23 -16 24 -12
rect 28 -16 29 -12
rect 23 -24 29 -16
rect 31 -24 32 -12
rect 36 -24 37 -12
rect 39 -24 40 -12
rect 44 -24 45 -12
rect 47 -24 48 -12
rect 63 -24 64 -12
rect 66 -24 67 -12
rect -51 -64 -48 -57
rect -46 -64 -45 -57
<< ndcontact >>
rect -48 -45 -44 -36
rect -40 -45 -36 -36
rect -53 -83 -49 -76
rect -45 -83 -41 -76
rect -27 -66 -23 -61
rect -13 -73 -9 -69
rect 0 -73 4 -61
rect 8 -73 12 -61
rect 16 -73 20 -61
rect 29 -73 33 -69
rect 42 -65 46 -61
rect 59 -51 63 -43
rect 67 -51 71 -43
<< pdcontact >>
rect -48 -24 -44 -12
rect -40 -24 -36 -12
rect -32 -24 -28 -12
rect -24 -24 -20 -12
rect -16 -24 -12 -12
rect -8 -16 -4 -12
rect 0 -24 4 -12
rect 8 -24 12 -12
rect 16 -24 20 -12
rect 24 -16 28 -12
rect 32 -24 36 -12
rect 40 -24 44 -12
rect 48 -24 52 -12
rect 59 -24 63 -12
rect 67 -24 71 -12
rect -55 -64 -51 -57
rect -45 -64 -41 -57
<< psubstratepcontact >>
rect -56 -44 -52 -40
<< nsubstratencontact >>
rect 78 -20 82 -16
rect -66 -67 -62 -63
<< polysilicon >>
rect -43 -12 -41 -10
rect -27 -12 -25 -10
rect -19 -12 -17 3
rect -11 -12 -9 -10
rect -3 -12 -1 12
rect 5 -12 7 12
rect 13 -12 15 12
rect 21 -12 23 12
rect 29 -12 31 -1
rect 37 -12 39 -10
rect 45 -12 47 -10
rect 64 -12 66 -10
rect -43 -28 -41 -24
rect -27 -26 -25 -24
rect -19 -26 -17 -24
rect -70 -30 -41 -28
rect -43 -36 -41 -30
rect -29 -28 -25 -26
rect -29 -45 -27 -28
rect -11 -32 -9 -24
rect -3 -41 -1 -24
rect -43 -48 -41 -45
rect -30 -47 -27 -45
rect -21 -43 -1 -41
rect -43 -50 -33 -48
rect -48 -57 -46 -55
rect -48 -69 -46 -64
rect -70 -71 -46 -69
rect -48 -76 -46 -71
rect -48 -90 -46 -83
rect -42 -90 -39 -86
rect -35 -91 -33 -50
rect -30 -75 -28 -47
rect -21 -61 -19 -43
rect 5 -46 7 -24
rect -3 -48 7 -46
rect 13 -46 15 -24
rect 21 -41 23 -24
rect 29 -26 31 -24
rect 37 -34 39 -24
rect 32 -36 39 -34
rect 21 -43 41 -41
rect 13 -48 23 -46
rect -16 -61 -14 -59
rect -8 -61 -6 -59
rect -3 -61 -1 -48
rect 5 -61 7 -59
rect 13 -61 15 -59
rect 21 -61 23 -48
rect 26 -59 27 -55
rect 26 -61 31 -59
rect 34 -61 36 -59
rect 39 -61 41 -43
rect 45 -45 47 -24
rect 64 -43 66 -24
rect 45 -47 52 -45
rect -21 -75 -19 -73
rect -16 -75 -14 -73
rect -30 -77 -27 -75
rect -29 -86 -27 -77
rect -8 -79 -6 -73
rect -3 -74 -1 -73
rect -3 -76 1 -74
rect -2 -78 1 -76
rect 5 -86 7 -73
rect -29 -88 7 -86
rect 13 -91 15 -73
rect 21 -80 23 -73
rect 26 -75 28 -73
rect 34 -86 36 -73
rect 39 -77 41 -73
rect 39 -79 46 -77
rect 44 -82 46 -79
rect 50 -91 52 -47
rect 64 -53 66 -51
rect -35 -93 52 -91
<< polycontact >>
rect -4 12 0 16
rect 4 12 8 16
rect 12 12 16 16
rect 20 12 24 16
rect -17 -1 -13 3
rect 28 -1 32 3
rect -74 -31 -70 -27
rect -33 -31 -29 -27
rect -12 -36 -8 -32
rect -74 -72 -70 -68
rect -46 -90 -42 -86
rect 28 -36 32 -32
rect -16 -59 -12 -55
rect 27 -59 31 -55
rect 60 -35 64 -31
rect -23 -79 -19 -75
rect -9 -83 -5 -79
rect -2 -82 2 -78
rect 20 -84 24 -80
rect 36 -86 40 -82
rect 43 -86 47 -82
rect -7 -109 -3 -105
rect 4 -107 8 -103
rect 12 -107 16 -103
rect 23 -109 27 -105
<< metal1 >>
rect -59 9 -56 16
rect -59 6 63 9
rect -48 -12 -44 6
rect -32 -4 -28 6
rect -13 -1 28 3
rect -32 -7 -4 -4
rect -32 -12 -28 -7
rect -8 -12 -4 -7
rect 24 -7 52 -4
rect 24 -12 28 -7
rect 48 -12 52 -7
rect -55 -24 -48 -12
rect -55 -40 -51 -24
rect -40 -27 -36 -24
rect -40 -31 -33 -27
rect -40 -36 -36 -31
rect -52 -44 -51 -40
rect -55 -57 -51 -44
rect -24 -43 -20 -24
rect -16 -26 -12 -24
rect 0 -26 4 -24
rect -16 -29 4 -26
rect 8 -43 12 -24
rect 16 -26 20 -24
rect 32 -26 36 -24
rect 16 -29 36 -26
rect 40 -43 44 -24
rect 59 -12 63 6
rect 74 7 78 16
rect 48 -31 52 -24
rect 67 -31 71 -24
rect 48 -35 60 -31
rect 67 -35 85 -31
rect -48 -48 -44 -45
rect -24 -46 44 -43
rect -48 -51 -31 -48
rect -66 -95 -62 -67
rect -59 -64 -55 -57
rect -59 -109 -56 -64
rect -45 -68 -41 -64
rect -45 -76 -41 -72
rect -53 -95 -49 -83
rect -35 -95 -31 -51
rect -27 -52 4 -49
rect -27 -61 -23 -52
rect 0 -61 4 -52
rect 16 -52 46 -49
rect 16 -61 20 -52
rect 42 -61 46 -52
rect -23 -105 -19 -79
rect -16 -76 -9 -73
rect -16 -95 -12 -76
rect -2 -95 2 -82
rect 20 -95 24 -84
rect -2 -99 8 -95
rect 4 -103 8 -99
rect -23 -109 -7 -105
rect 12 -99 24 -95
rect 29 -95 33 -73
rect 49 -74 52 -35
rect 67 -43 71 -35
rect 43 -77 52 -74
rect 12 -103 16 -99
rect 43 -105 47 -86
rect 59 -95 63 -51
rect 27 -109 47 -105
rect 74 -109 78 -99
<< m2contact >>
rect 32 -1 36 3
rect -78 -31 -74 -27
rect -12 -40 -8 -36
rect 28 -40 32 -36
rect 74 3 78 7
rect 74 -20 78 -16
rect -78 -72 -74 -68
rect -66 -99 -62 -95
rect -45 -72 -41 -68
rect -42 -90 -38 -86
rect -53 -99 -49 -95
rect -20 -59 -16 -55
rect -12 -59 -8 -55
rect 23 -59 27 -55
rect -35 -99 -31 -95
rect 8 -77 12 -73
rect -9 -87 -5 -83
rect -16 -99 -12 -95
rect 39 -78 43 -74
rect 36 -90 40 -86
rect 29 -99 33 -95
rect 59 -99 63 -95
rect 74 -99 78 -95
<< metal2 >>
rect 36 -1 56 3
rect -12 -55 -8 -40
rect 28 -52 32 -40
rect 23 -55 32 -52
rect -31 -59 -20 -55
rect -16 -59 -12 -55
rect -8 -58 23 -55
rect -8 -59 5 -58
rect 15 -59 23 -58
rect 27 -59 32 -55
rect -31 -68 -28 -59
rect -41 -72 -28 -68
rect 12 -77 39 -74
rect -9 -83 -5 -79
rect -2 -82 2 -78
rect -43 -90 -42 -87
rect -38 -87 -9 -86
rect 53 -86 56 -1
rect 74 -16 78 3
rect 59 -51 63 -43
rect 67 -51 71 -43
rect -5 -87 18 -86
rect 26 -87 36 -86
rect -38 -90 36 -87
rect 40 -90 56 -86
rect 74 -95 78 -20
rect -62 -99 -53 -95
rect -49 -99 -35 -95
rect -31 -99 -16 -95
rect -12 -99 29 -95
rect 33 -99 59 -95
rect 63 -99 74 -95
<< m3contact >>
rect -82 -31 -78 -27
rect -82 -72 -78 -68
<< metal3 >>
rect -83 -27 -77 -26
rect -83 -31 -82 -27
rect -78 -31 -77 -27
rect -83 -32 -77 -31
rect -83 -68 -77 -67
rect -83 -72 -82 -68
rect -78 -72 -77 -68
rect -83 -73 -77 -72
<< labels >>
rlabel metal1 50 -35 50 -35 1 _f
rlabel polysilicon -60 -29 -60 -29 1 a
rlabel polysilicon 30 -3 30 -3 1 t1
rlabel metal1 73 -33 73 -33 7 f
rlabel polysilicon -60 -70 -60 -70 3 b
rlabel polycontact -2 14 -2 14 1 g1
rlabel polycontact 6 14 6 14 1 g2
rlabel polycontact 14 14 14 14 1 g3
rlabel polycontact 22 14 22 14 1 g4
rlabel metal1 -59 12 -56 16 1 Vdd!
rlabel metal1 74 12 78 16 1 GND!
rlabel metal1 81 -35 85 -31 7 f
<< end >>
